// Define your enumerated type(s) here

class yapp_packet extends uvm_sequence_item;

// Define the protocol data

// Define control knobs

// Enable automation of the packet's fields

// Define packet constraints

// Add methods for parity calculation and class construction

endclass: yapp_packet
