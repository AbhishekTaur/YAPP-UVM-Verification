/*-----------------------------------------------------------------
File name     : hbus_pkg.sv
Developers    : Kathleen Meade
Created       : Wed Mar 11 2009
Description   :
Notes         :
-------------------------------------------------------------------
Copyright 2009 (c) Cadence Design Systems
-----------------------------------------------------------------*/

`ifndef HBUS_PKG_SV
`define HBUS_PKG_SV

package hbus_pkg;

 import uvm_pkg::*;
 `include "uvm_macros.svh"

 `include "hbus.svh"

endpackage : hbus_pkg

`endif // HBUS_PKG_SV
