/*-----------------------------------------------------------------
File name     : channel_pkg.sv
Developers    : Kathleen Meade
Created       : March 11, 2009
Description   : This creates a package for the channel OVC
Notes         :
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2009 
-----------------------------------------------------------------*/

package channel_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "channel.svh"

endpackage : channel_pkg
