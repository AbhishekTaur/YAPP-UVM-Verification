/*-----------------------------------------------------------------
File name     : yapp_pkt_pkg.sv
Developers    : Kathleen Meade
Created       : March 11, 2009
Description   : This creates a package for the YAPP packet
Notes         :
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2009 
-----------------------------------------------------------------*/

package yapp_pkt_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "yapp_packet.sv"

endpackage : yapp_pkt_pkg
