/*-----------------------------------------------------------------
File name     : yapp.svh
Developers    : Brian Dickinson
Created       : 01/06/09
Description   : This file imports all the files of the simple YAPP OVC.
Notes         :
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2009
-----------------------------------------------------------------*/

`include "yapp_packet.sv"
`include "yapp_tx_monitor.sv"
`include "yapp_tx_sequencer.sv"
`include "yapp_tx_seqs.sv"
`include "yapp_tx_driver.sv"
`include "yapp_tx_agent.sv"
`include "yapp_env.sv"

