// CDNS GIT SHA "UVM_1_1-78-g07f7862" last-MERGED-state from Accellera "UVM-1.0p1-5-g16015a6" 
