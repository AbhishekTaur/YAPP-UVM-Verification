/*-------------------------------------------------------------------------
File name   : router.svh
Title       : Module UVC Files
----------------------------------------------------------------------*/

import yapp_pkt_pkg::*;
// import HBUS package for visibility of HBUS data item
import hbus_pkg::*;
`include "router_scoreboard.sv"
`include "router_reference.sv"
`include "router_module_env.sv"
