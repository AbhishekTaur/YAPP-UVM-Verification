/*-----------------------------------------------------------------
File name     : router_module_pkg.sv
Developers    : Abhishek Taur
Created       : 06/14/19
Description   : Package includes router module UVC files
Notes         :
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2011
-----------------------------------------------------------------*/
package router_module_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "router_module.svh"

endpackage

