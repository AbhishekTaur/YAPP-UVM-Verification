/*-----------------------------------------------------------------
File name     : yapp_pkg.sv
Developers    : Brian Dickinson
Created       : 01/04/11
Description   : Package includes YAPP UVC header file
Notes         :
-------------------------------------------------------------------
Copyright Cadence Design Systems (c)2011
-----------------------------------------------------------------*/
package yapp_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "yapp.svh"

endpackage
