module packet_test;
  import packet_classes::*;

  // step 1:
  // construct, load and print a basic packet instance


  // step 2:
  // create an array of base class  
  // create handles for every packet type
  // randomly assign packet sub-class instances to base array elements
  //   use randomize and assignment to set packet data
  // print  array

endmodule
   

